// PLL.v

// Generated using ACDS version 13.0 156 at 2018.06.04.20:03:36

`timescale 1 ps / 1 ps
module PLL (
		input  wire  clk_in_clk,  // clk_in.clk
		input  wire  reset_reset, //  reset.reset
		output wire  c0_clk,      //     c0.clk
		output wire  clk_c1_clk   // clk_c1.clk
	);

	PLL_altpll_0 altpll_0 (
		.clk       (clk_in_clk),  //       inclk_interface.clk
		.reset     (reset_reset), // inclk_interface_reset.reset
		.read      (),            //             pll_slave.read
		.write     (),            //                      .write
		.address   (),            //                      .address
		.readdata  (),            //                      .readdata
		.writedata (),            //                      .writedata
		.c0        (c0_clk),      //                    c0.clk
		.c1        (clk_c1_clk),  //                    c1.clk
		.areset    (),            //        areset_conduit.export
		.locked    (),            //        locked_conduit.export
		.phasedone ()             //     phasedone_conduit.export
	);

endmodule
